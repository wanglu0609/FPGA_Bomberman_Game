module bird_sprite(output logic [9:0] rgb[0:31][0:31]);
assign rgb = '{
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd1,9'd2,9'd1,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd3,9'd4,9'd5,9'd6,9'd7,9'd8,9'd9,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd10,9'd10,9'd11,9'd12,9'd0,9'd0,9'd0,9'd0,9'd0,9'd8,9'd4,9'd13,9'd14,9'd15,9'd16,9'd17,9'd6,9'd6,9'd5,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd18,9'd19,9'd18,9'd20,9'd21,9'd21,9'd22,9'd21,9'd12,9'd23,9'd5,9'd24,9'd25,9'd26,9'd27,9'd28,9'd29,9'd30,9'd31,9'd32,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd33,9'd34,9'd24,9'd24,9'd35,9'd36,9'd37,9'd11,9'd12,9'd12,9'd38,9'd39,9'd40,9'd41,9'd26,9'd26,9'd26,9'd42,9'd43,9'd44,9'd45,9'd46,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd18,9'd11,9'd47,9'd37,9'd34,9'd34,9'd36,9'd48,9'd37,9'd11,9'd12,9'd49,9'd39,9'd50,9'd27,9'd26,9'd26,9'd26,9'd51,9'd52,9'd44,9'd9,9'd5,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd34,9'd22,9'd22,9'd22,9'd22,9'd11,9'd53,9'd54,9'd53,9'd37,9'd12,9'd12,9'd5,9'd4,9'd55,9'd26,9'd26,9'd26,9'd26,9'd28,9'd27,9'd51,9'd56,9'd57,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd19,9'd58,9'd58,9'd22,9'd59,9'd60,9'd61,9'd62,9'd53,9'd63,9'd48,9'd64,9'd65,9'd5,9'd24,9'd29,9'd26,9'd26,9'd26,9'd26,9'd28,9'd26,9'd66,9'd43,9'd67,9'd68,9'd69,9'd0
},
'{
9'd0,9'd0,9'd0,9'd35,9'd22,9'd58,9'd59,9'd70,9'd71,9'd72,9'd73,9'd72,9'd71,9'd74,9'd53,9'd53,9'd75,9'd5,9'd16,9'd41,9'd26,9'd26,9'd26,9'd26,9'd26,9'd28,9'd76,9'd43,9'd77,9'd78,9'd5,9'd0
},
'{
9'd0,9'd0,9'd79,9'd58,9'd58,9'd80,9'd22,9'd81,9'd82,9'd83,9'd84,9'd83,9'd85,9'd86,9'd87,9'd54,9'd88,9'd6,9'd15,9'd26,9'd26,9'd26,9'd26,9'd26,9'd28,9'd26,9'd43,9'd43,9'd56,9'd6,9'd6,9'd0
},
'{
9'd0,9'd89,9'd35,9'd21,9'd12,9'd80,9'd22,9'd90,9'd91,9'd92,9'd93,9'd93,9'd84,9'd94,9'd95,9'd96,9'd9,9'd7,9'd97,9'd26,9'd26,9'd26,9'd26,9'd26,9'd27,9'd98,9'd43,9'd44,9'd99,9'd39,9'd88,9'd0
},
'{
9'd0,9'd79,9'd20,9'd12,9'd11,9'd12,9'd58,9'd100,9'd101,9'd102,9'd103,9'd104,9'd93,9'd83,9'd85,9'd95,9'd105,9'd106,9'd97,9'd27,9'd28,9'd26,9'd27,9'd26,9'd28,9'd107,9'd43,9'd52,9'd108,9'd39,9'd65,9'd0
},
'{
9'd0,9'd109,9'd47,9'd20,9'd110,9'd70,9'd58,9'd111,9'd112,9'd113,9'd114,9'd115,9'd116,9'd117,9'd118,9'd111,9'd119,9'd120,9'd109,9'd121,9'd14,9'd26,9'd122,9'd27,9'd28,9'd76,9'd43,9'd123,9'd124,9'd39,9'd64,9'd0
},
'{
9'd47,9'd4,9'd37,9'd80,9'd53,9'd70,9'd59,9'd125,9'd126,9'd127,9'd128,9'd129,9'd130,9'd131,9'd132,9'd133,9'd134,9'd135,9'd78,9'd24,9'd28,9'd27,9'd107,9'd52,9'd136,9'd137,9'd138,9'd139,9'd6,9'd9,9'd10,9'd0
},
'{
9'd37,9'd24,9'd75,9'd48,9'd53,9'd140,9'd74,9'd141,9'd142,9'd127,9'd113,9'd128,9'd143,9'd143,9'd144,9'd141,9'd145,9'd129,9'd146,9'd135,9'd147,9'd41,9'd148,9'd43,9'd123,9'd78,9'd149,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd47,9'd121,9'd17,9'd35,9'd53,9'd48,9'd74,9'd150,9'd132,9'd126,9'd127,9'd151,9'd152,9'd126,9'd153,9'd154,9'd155,9'd156,9'd157,9'd131,9'd149,9'd124,9'd31,9'd158,9'd139,9'd124,9'd68,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd70,9'd79,9'd40,9'd24,9'd54,9'd159,9'd60,9'd160,9'd161,9'd162,9'd156,9'd163,9'd164,9'd102,9'd165,9'd166,9'd163,9'd167,9'd156,9'd168,9'd4,9'd5,9'd9,9'd124,9'd169,9'd170,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd80,9'd23,9'd40,9'd5,9'd17,9'd17,9'd17,9'd62,9'd171,9'd162,9'd172,9'd156,9'd173,9'd174,9'd175,9'd128,9'd163,9'd156,9'd172,9'd126,9'd176,9'd177,9'd178,9'd32,9'd117,9'd86,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd140,9'd18,9'd4,9'd40,9'd4,9'd63,9'd17,9'd159,9'd179,9'd154,9'd151,9'd114,9'd157,9'd180,9'd181,9'd115,9'd182,9'd114,9'd173,9'd174,9'd183,9'd184,9'd180,9'd92,9'd185,9'd186,9'd187,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd11,9'd121,9'd124,9'd4,9'd188,9'd63,9'd159,9'd189,9'd190,9'd191,9'd192,9'd180,9'd193,9'd192,9'd115,9'd194,9'd194,9'd195,9'd196,9'd197,9'd198,9'd193,9'd199,9'd200,9'd85,9'd187,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd21,9'd36,9'd121,9'd108,9'd69,9'd201,9'd202,9'd189,9'd160,9'd203,9'd103,9'd155,9'd102,9'd126,9'd173,9'd194,9'd157,9'd204,9'd155,9'd205,9'd205,9'd206,9'd129,9'd145,9'd207,9'd208,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd47,9'd11,9'd36,9'd75,9'd5,9'd209,9'd54,9'd140,9'd210,9'd82,9'd211,9'd166,9'd212,9'd213,9'd126,9'd173,9'd214,9'd215,9'd216,9'd152,9'd216,9'd217,9'd164,9'd218,9'd185,9'd187,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd58,9'd36,9'd65,9'd75,9'd17,9'd159,9'd60,9'd219,9'd219,9'd220,9'd221,9'd156,9'd213,9'd173,9'd167,9'd222,9'd165,9'd223,9'd224,9'd225,9'd226,9'd222,9'd129,9'd227,9'd96,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd22,9'd37,9'd65,9'd140,9'd17,9'd60,9'd60,9'd219,9'd228,9'd229,9'd167,9'd126,9'd114,9'd166,9'd230,9'd231,9'd232,9'd233,9'd234,9'd226,9'd130,9'd129,9'd183,9'd235,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd110,9'd12,9'd110,9'd70,9'd140,9'd189,9'd74,9'd74,9'd179,9'd133,9'd151,9'd163,9'd174,9'd173,9'd191,9'd236,9'd237,9'd238,9'd237,9'd239,9'd157,9'd126,9'd227,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd47,9'd58,9'd11,9'd70,9'd70,9'd59,9'd240,9'd219,9'd72,9'd191,9'd241,9'd214,9'd200,9'd197,9'd242,9'd243,9'd244,9'd239,9'd241,9'd245,9'd128,9'd203,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd58,9'd12,9'd58,9'd58,9'd12,9'd22,9'd74,9'd22,9'd86,9'd184,9'd184,9'd101,9'd112,9'd128,9'd246,9'd164,9'd218,9'd182,9'd157,9'd229,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd11,9'd22,9'd22,9'd22,9'd58,9'd22,9'd74,9'd247,9'd80,9'd248,9'd249,9'd250,9'd249,9'd249,9'd251,9'd252,9'd252,9'd251,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd47,9'd22,9'd58,9'd22,9'd58,9'd58,9'd22,9'd247,9'd247,9'd247,9'd253,9'd48,9'd211,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd11,9'd22,9'd22,9'd22,9'd22,9'd140,9'd11,9'd22,9'd247,9'd22,9'd22,9'd22,9'd22,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd58,9'd22,9'd22,9'd80,9'd36,9'd11,9'd22,9'd58,9'd12,9'd12,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd12,9'd12,9'd0,9'd0,9'd47,9'd47,9'd47,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
}};
endmodule
