module  Color_Mapper_Final (
	input [9:0] Avatar_X_1, Avatar_Y_1, Avatar_Step_1,     // Ball coordinates
	            Avatar_X_2, Avatar_Y_2, Avatar_Step_2,
					Draw_X, Draw_Y,      // Coordinates of current drawing pixel
	input [1:0] Avatar_Dir_1,  Avatar_Dir_2, state,
   input [143:0] Wall_Map, Tree_Map, Treasure_Map, Bomb_Map, Flame_Map,
	input [7:0] score_0, score_1,
	input Player_choose, Winner,
	output logic [7:0] VGA_R, VGA_G, VGA_B // VGA RGB output
);
 
	logic [7:0] c_table[0:33][0:2];
	logic [7:0] Red, Green, Blue;
	logic [7:0] av_index_1, av_index_2, temp_1, temp_2,
	            tile_index, small_index, big_index;
	logic [7:0] avf [0:179][0:39];
   logic [7:0] avr [0:179][0:39];
	logic [7:0] avb [0:179][0:39];
	logic [7:0] ground [0:39][0:39];
	logic [7:0] tree [0:39][0:39];
	logic [7:0] bomb_1 [0:27][0:27];
	logic [7:0] flame_1 [0:27][0:27];
	logic [7:0] wall [0:39][0:39];
	logic front_on_2, right_on_2, left_on_2, back_on_2, wall_on, tree_on, flame_on, bomb_on, again_on,
	      front_on_1, right_on_1, left_on_1, back_on_1, av_1, av_2, coin_on, player1_on, player2_on, final_on;
   logic [3:0] score_on;
   logic [10:0] sprite_addr;
   logic [7:0] sprite_data;
	logic [5:0] addr_scene;
	logic [3:0] addr_2;
	logic [97:0] sprite_scene,sprite_2;
	
	
   font_rom newfont(.addr(sprite_addr), .data(sprite_data));	
	big_font newscene(.addr(addr_scene), .data(sprite_scene));
   again_font again_1(.addr(addr_2), .data(sprite_2));	

	color_table color(.colors(c_table));
	front ava_f(.index(avf));
	right ava_r(.index(avr));
	back ava_b(.index(avb));
	tile background(.index(ground));
	Solid solidwall(.index(wall));
	flame fire(.index(flame_1));
	bomb_sprites explode(.index(bomb_1));
	exploded EB(.index(tree));

	int Char_X_1, Char_Y_1, loc_x_1, loc_y_1, Char_X_2, Char_Y_2, loc_x_2, loc_y_2, move_1, move_2;
	int step_1, step_2, t1, t2, width, height, cell_x, cell_y;
	int score_index_0, score_index_1, score_x_0, score_x_1;
	int player_x, player_1_y, player_2_y, win_x, win_y, again_x, again_y;
	assign Char_X_1 = Avatar_X_1;
	assign Char_Y_1 = Avatar_Y_1;
   assign Char_X_2 = Avatar_X_2;
	assign Char_Y_2 = Avatar_Y_2;
	assign width = 20;
	assign height = 40;
	assign loc_x_1 = Draw_X - Char_X_1 + width;
	assign loc_y_1 = Draw_Y - Char_Y_1 + height;
   assign loc_x_2 = Draw_X - Char_X_2 + width;
	assign loc_y_2 = Draw_Y - Char_Y_2 + height;
	assign step_1 = Avatar_Step_1;
	assign step_2 = Avatar_Step_2;
	assign move_1 = (step_1/4) % 2;
	assign move_2 = (step_2/4) % 2;
	assign t1 = Draw_X % 40;
   assign t2 = Draw_Y % 40;
	assign cell_x = Draw_X / 40;
	assign cell_y = Draw_Y / 40;
	assign score_index_0 = Draw_Y - 212;
	assign score_index_1 = Draw_Y - 252;
	assign score_x_0 = Draw_X - 596;
	assign score_x_1 = Draw_X - 611;
	assign player_x = Draw_X - 271;
   assign player_1_y = Draw_Y - 192;
   assign player_2_y = Draw_Y - 272;
	assign win_x = Draw_X - 222;
	assign win_y = Draw_Y - 224;
	assign again_x = Draw_X - 271;
	assign again_y = Draw_Y - 280;
	
	assign tile_index = ground[t2][t1];
	
	assign VGA_R = Red;
	assign VGA_G = Green;
	assign VGA_B = Blue;

	

	always_comb
	begin : find_index

		if(state == 2'b01 && Draw_X >= Char_X_1 - width && Draw_X < Char_X_1 + width && Draw_Y >= Char_Y_1 - height && Draw_Y < Char_Y_1 + width) 
		begin
			if(Avatar_Dir_1==2'b00)
			begin 
			   front_on_1 = 1'b1;
			   av_1 = 1'b1; 
	         right_on_1= 1'b0; 
	         left_on_1= 1'b0; 
	         back_on_1= 1'b0; 
				
			end
			else if(Avatar_Dir_1==2'b01)
			begin 
			   back_on_1 = 1'b1;
			   av_1 = 1'b1;
	         front_on_1= 1'b0; 
	         right_on_1= 1'b0; 
	         left_on_1= 1'b0; 
			end
			else if(Avatar_Dir_1==2'b10)
			begin 
			   left_on_1 = 1'b1;
			   av_1 = 1'b1;
	         front_on_1= 1'b0; 
	         right_on_1= 1'b0; 
	         back_on_1= 1'b0; 
			end
			else
			begin 
			   right_on_1 = 1'b1;
			   av_1 = 1'b1;
	         front_on_1= 1'b0; 
	         left_on_1= 1'b0; 
	         back_on_1= 1'b0; 
			end

		end
		else
		begin
		   av_1 = 1'b0;
	      front_on_1= 1'b0; 
       	right_on_1= 1'b0; 
	      left_on_1= 1'b0; 
	      back_on_1= 1'b0; 
		end
		
		if(state == 2'b01 && Draw_X >= Char_X_2 - width && Draw_X < Char_X_2 + width && Draw_Y >= Char_Y_2 - height && Draw_Y < Char_Y_2 + width) 
		begin
		   if(Avatar_Dir_2==2'b00)
			begin 
			   front_on_2 = 1'b1;
			   av_2 = 1'b1;
	         right_on_2 = 1'b0; 
	         left_on_2 =  1'b0;
	         back_on_2 = 1'b0;
			end
			else if(Avatar_Dir_2==2'b01)
			begin 
			   back_on_2 = 1'b1;
			   av_2 = 1'b1;
				front_on_2 = 1'b0;
	         right_on_2 = 1'b0; 
	         left_on_2 =  1'b0;
			end
			else if(Avatar_Dir_2==2'b10)
			begin 
			   left_on_2 = 1'b1;
			   av_2 = 1'b1;
				front_on_2 = 1'b0;
	         right_on_2 = 1'b0; 
         	back_on_2 = 1'b0;
			end
			else
			begin 
			   right_on_2 = 1'b1;
			   av_2 = 1'b1;
				front_on_2 = 1'b0;
				left_on_2 =  1'b0;
				back_on_2 = 1'b0;
			end

		end
		else
		begin
		   av_2 = 1'b0;
		   left_on_2 = 1'b0;
			front_on_2 = 1'b0;
	      right_on_2 = 1'b0; 
         back_on_2 = 1'b0;
		end
		
		if((state == 2'b01) && (Draw_X < 480)&&(Bomb_Map[cell_y*12+cell_x]))
		begin
		   bomb_on = 1'b1;
			wall_on = 1'b0;
			tree_on = 1'b0;
			flame_on = 1'b0;
			coin_on = 1'b0;
		end
		else if((state == 2'b01) && (Draw_X < 480)&&(Wall_Map[cell_y*12+cell_x]))
		begin
		   wall_on = 1'b1;
			bomb_on = 1'b0;
			tree_on = 1'b0;
			flame_on = 1'b0;
			coin_on = 1'b0;
		end
		else if((state == 2'b01) && (Draw_X < 480)&&(Flame_Map[cell_y*12+cell_x]))
		begin
		   flame_on = 1'b1;
			bomb_on = 1'b0;
			wall_on = 1'b0;
			tree_on = 1'b0;
			coin_on = 1'b0;
		end
		else if((state == 2'b01) && (Draw_X < 480)&&(Tree_Map[cell_y*12+cell_x]))
		begin
		   tree_on = 1'b1;
			bomb_on = 1'b0;
			wall_on = 1'b0;
			flame_on = 1'b0;
			coin_on = 1'b0;
		end
		else if((state == 2'b01) && (Draw_X<480)&&(Treasure_Map[cell_y*12+cell_x])&&(Draw_X>cell_x*40+12)&&(Draw_X<=cell_x*40+28)&&(Draw_Y>cell_y*40+12)&&(Draw_Y<=cell_y*40+28))
		begin
		   coin_on = 1'b1;
		   tree_on = 1'b0;
			bomb_on = 1'b0;
			wall_on = 1'b0;
			flame_on = 1'b0;
		end
		else 
		begin
			coin_on = 1'b0;
			bomb_on = 1'b0;
			wall_on = 1'b0;
			tree_on = 1'b0;
			flame_on = 1'b0;
		end
		if(state == 2'b01 && Draw_X > 596 && Draw_X <= 604 && Draw_Y > 212 && Draw_Y < 228)
		   score_on = 4'b0010;
		else if(state == 2'b01 && Draw_X > 611 && Draw_X <= 619 && Draw_Y > 212 && Draw_Y <= 228)
		   score_on = 4'b0001;	
		else if(state == 2'b01 && Draw_X > 596 && Draw_X <= 604 && Draw_Y > 252 && Draw_Y <= 268)
		   score_on = 4'b1000;
		else if(state == 2'b01 && Draw_X > 611 && Draw_X <= 619 && Draw_Y > 252 && Draw_Y <= 268)
		   score_on = 4'b0100;
		else
		   score_on = 4'b0000;
			
		if(state == 2'b00)
		begin
		   if(Draw_X > 271 && Draw_X <= 369 && Draw_Y > 192 && Draw_Y <= 208)
			begin
		      player1_on = 1'b1;
				player2_on = 1'b0;
			   final_on = 1'b0;
				again_on = 1'b0;
			end
			else if(Draw_X > 271 && Draw_X <= 369 && Draw_Y > 272 && Draw_Y <= 288)
			begin
		      player1_on = 1'b0;
				player2_on = 1'b1;
			   final_on = 1'b0;
				again_on = 1'b0;
			end
			else
			begin
		      player1_on = 1'b0;
				player2_on = 1'b0;
			   final_on = 1'b0;
				again_on = 1'b0;
			end
		end
		else if(state == 2'b01)
		begin
		   player1_on = 1'b0;
			player2_on = 1'b0;
			final_on = 1'b0;
			again_on = 1'b0;
		end
		else if(state == 2'b10)
		begin
		   if(Draw_X > 271 && Draw_X <= 369 && Draw_Y > 280 && Draw_Y <= 296)
			begin
		      player1_on = 1'b0;
			   player2_on = 1'b0;
			   final_on = 1'b0;
				again_on = 1'b1;
			end
		   else if(Draw_X > 222 && Draw_X <= 418 && Draw_Y > 224 && Draw_Y <= 256)
			begin
		      player1_on = 1'b0;
			   player2_on = 1'b0;
			   final_on = 1'b1;
				again_on = 1'b0;
			end
			else
			begin
		      player1_on = 1'b0;
			   player2_on = 1'b0;
			   final_on = 1'b0;
				again_on = 1'b0;
			end
		end
		else
		begin
		   player1_on = 1'b0;
			player2_on = 1'b0;
			final_on = 1'b0;
			again_on = 1'b0;
		end
	end

	
	
	

	always_comb
   begin : color_picker
	   if (front_on_1 == 1'b1) 
		begin
		   if((step_1<2)||(step_1>37))
		   begin
			    av_index_1 = avf[loc_y_1+60][loc_x_1];
		   end
	   	else if (move_1 == 0)
		   begin
             av_index_1 = avf[loc_y_1+120][loc_x_1];
			end
	   	else
		   begin
             av_index_1 = avf[loc_y_1][loc_x_1];
			end
			
		end
		else if (back_on_1 == 1'b1) 
		begin
		   if((step_1<2)||(step_1>37))
		   begin
			    av_index_1 = avb[loc_y_1+60][loc_x_1];
		   end
	   	else if (move_1 == 0)
		   begin
             av_index_1 = avb[loc_y_1+120][loc_x_1];
			end
	   	else
		   begin
             av_index_1 = avb[loc_y_1][loc_x_1];
			end
			
		end
		else if (right_on_1 == 1'b1) 
		begin
		   if((step_1<2)||(step_1>37))
		   begin
			    av_index_1 = avr[loc_y_1+60][loc_x_1];
		   end
	   	else if (move_1 == 0)
		   begin
             av_index_1 = avr[loc_y_1+120][loc_x_1];
			end
	   	else
		   begin
             av_index_1 = avr[loc_y_1][loc_x_1];
			end
			
		end
		else if (left_on_1 == 1'b1) 
		begin
		   if((step_1<2)||(step_1>37))
		   begin
			    av_index_1 = avr[loc_y_1+60][39-loc_x_1];
		   end
	   	else if (move_1 == 0)
		   begin
             av_index_1 = avr[loc_y_1+120][39-loc_x_1];
			end
	   	else
		   begin
             av_index_1 = avr[loc_y_1][39-loc_x_1];
			end
			
		end
		else
		begin
		   av_index_1 = 0;
		end
	   if (front_on_2 == 1'b1) 
		begin
		   if((step_2<2)||(step_2>37))
		   begin
			    av_index_2 = avf[loc_y_2+60][loc_x_2];
		   end
	   	else if (move_2 == 0)
		   begin
             av_index_2 = avf[loc_y_2+120][loc_x_2];
			end
	   	else
		   begin
             av_index_2 = avf[loc_y_2][loc_x_2];
			end
			
		end
		else if (back_on_2 == 1'b1) 
		begin
		   if((step_2<2)||(step_2>37))
		   begin
			    av_index_2 = avb[loc_y_2+60][loc_x_2];
		   end
	   	else if (move_2 == 0)
		   begin
             av_index_2 = avb[loc_y_2+120][loc_x_2];
			end
	   	else
		   begin
             av_index_2 = avb[loc_y_2][loc_x_2];
			end
			
		end
		else if (right_on_2 == 1'b1) 
		begin
		   if((step_2<2)||(step_2>37))
		   begin
			    av_index_2 = avr[loc_y_2+60][loc_x_2];
		   end
	   	else if (move_2 == 0)
		   begin
             av_index_2 = avr[loc_y_2+120][loc_x_2];
			end
	   	else
		   begin
             av_index_2 = avr[loc_y_2][loc_x_2];
			end
			
		end
		else if (left_on_2 == 1'b1) 
		begin
		   if((step_2<2)||(step_2>37))
		   begin
			    av_index_2 = avr[loc_y_2+60][39-loc_x_2];
		   end
	   	else if (move_2 == 0)
		   begin
             av_index_2 = avr[loc_y_2+120][39-loc_x_2];
			end
	   	else
		   begin
             av_index_2 = avr[loc_y_2][39-loc_x_2];
			end
			
		end
		else
		begin
		   av_index_2 = 0;
		end		
			
		if(bomb_on == 1'b1)
		begin
			small_index =  bomb_1[t2-6][t1-6];
			big_index = 0;
		end
		else if(tree_on == 1'b1)
		begin
			big_index =  tree[t2][t1];
			small_index = 0;
		end
		else if(wall_on == 1'b1)
		begin
		   big_index = wall[t2][t1];
			small_index = 0;
		end
		else if(flame_on == 1'b1)
		begin
		   small_index = flame_1[t2-6][t1-6];
			big_index = 0;
		end
		else
		begin
			big_index = 0;
			small_index = 0;
		end
		
		
		if(score_on[0])
		begin
		    case(score_0%10)
		    4'd0: begin
            sprite_addr = score_index_0 + 16* 'h30;
          end		   
			 4'd1: begin
            sprite_addr = score_index_0 + 16* 'h31;
          end
			 4'd2: begin
            sprite_addr = score_index_0 + 16* 'h32;
          end
			 4'd3: begin
            sprite_addr = score_index_0 + 16* 'h33;
          end
			 4'd4: begin
            sprite_addr = score_index_0 + 16* 'h34;
          end
			 4'd5: begin
            sprite_addr = score_index_0 + 16* 'h35;
          end
			 4'd6: begin
            sprite_addr = score_index_0 + 16* 'h36;
          end
			 4'd7: begin
            sprite_addr = score_index_0 + 16* 'h37;
          end
			 4'd8: begin
            sprite_addr = score_index_0 + 16* 'h38;
          end
			 4'd9: begin
            sprite_addr = score_index_0 + 16* 'h39;
          end
			 default:
			   sprite_addr = 0;
		    endcase
		end
		else if(score_on[1])
		begin
		    case((score_0/10)%10)
		    4'd0: begin
            sprite_addr = score_index_0 + 16* 'h30;
          end		   
			 4'd1: begin
            sprite_addr = score_index_0 + 16* 'h31;
          end
			 4'd2: begin
            sprite_addr = score_index_0 + 16* 'h32;
          end
			 4'd3: begin
            sprite_addr = score_index_0 + 16* 'h33;
          end
			 4'd4: begin
            sprite_addr = score_index_0 + 16* 'h34;
          end
			 4'd5: begin
            sprite_addr = score_index_0 + 16* 'h35;
          end
			 4'd6: begin
            sprite_addr = score_index_0 + 16* 'h36;
          end
			 4'd7: begin
            sprite_addr = score_index_0 + 16* 'h37;
          end
			 4'd8: begin
            sprite_addr = score_index_0 + 16* 'h38;
          end
			 4'd9: begin
            sprite_addr = score_index_0 + 16* 'h39;
          end
			 default:
			   sprite_addr = 0;
		    endcase
		end
		else if(score_on[2])
		begin
		    case(score_1%10)
		    4'd0: begin
            sprite_addr = score_index_1 + 16* 'h30;
          end		   
			 4'd1: begin
            sprite_addr = score_index_1 + 16* 'h31;
          end
			 4'd2: begin
            sprite_addr = score_index_1 + 16* 'h32;
          end
			 4'd3: begin
            sprite_addr = score_index_1 + 16* 'h33;
          end
			 4'd4: begin
            sprite_addr = score_index_1 + 16* 'h34;
          end
			 4'd5: begin
            sprite_addr = score_index_1 + 16* 'h35;
          end
			 4'd6: begin
            sprite_addr = score_index_1 + 16* 'h36;
          end
			 4'd7: begin
            sprite_addr = score_index_1 + 16* 'h37;
          end
			 4'd8: begin
            sprite_addr = score_index_1 + 16* 'h38;
          end
			 4'd9: begin
            sprite_addr = score_index_1 + 16* 'h39;
          end
			 default:
			   sprite_addr = 0;
		    endcase
		end
		else if(score_on[3])
		begin
		    case((score_1/10)%10)
		    4'd0: begin
            sprite_addr = score_index_1 + 16* 'h30;
          end		   
			 4'd1: begin
            sprite_addr = score_index_1 + 16* 'h31;
          end
			 4'd2: begin
            sprite_addr = score_index_1 + 16* 'h32;
          end
			 4'd3: begin
            sprite_addr = score_index_1 + 16* 'h33;
          end
			 4'd4: begin
            sprite_addr = score_index_1 + 16* 'h34;
          end
			 4'd5: begin
            sprite_addr = score_index_1 + 16* 'h35;
          end
			 4'd6: begin
            sprite_addr = score_index_1 + 16* 'h36;
          end
			 4'd7: begin
            sprite_addr = score_index_1 + 16* 'h37;
          end
			 4'd8: begin
            sprite_addr = score_index_1 + 16* 'h38;
          end
			 4'd9: begin
            sprite_addr = score_index_1 + 16* 'h39;
          end
			 default:
			   sprite_addr = 0;
		    endcase
		end
		else if(coin_on)
		begin
		    sprite_addr = t2 - 12 + 16* 'h24;
		end
		else
		    sprite_addr = 0;
		if(player1_on)
		    addr_scene = player_1_y + 32;
		else if(player2_on)
		    addr_scene = player_2_y + 48;
		else if((final_on == 1'b1) && (Winner == 1'b0))
		    addr_scene = win_y/2; 
		else if((final_on == 1'b1)&&(Winner == 1'b1))
		    addr_scene = win_y/2  + 16;
		else
		    addr_scene = 0;
		if((again_on == 1'b1))
		    addr_2 = Draw_Y - 280;
		else addr_2 = 0;
	end 

	



	always_comb
	begin : RGB_Display
		if ((av_1 == 1'b1) && (av_index_1 != 0)) 
		begin
			Red = c_table[av_index_1][0];
			Green = c_table[av_index_1][1];
			Blue = c_table[av_index_1][2];
		end
		else if((av_2 == 1'b1) && (av_index_2 != 0)) 
		begin
		   if(av_index_2 == 8'd3)
			begin
			   Red = 8'd51;
			   Green = 8'd255;
			   Blue = 8'd255;
			end
			else
			begin
			   Red = c_table[av_index_2][0];
			   Green = c_table[av_index_2][1];
			   Blue = c_table[av_index_2][2];
			end
		end
		else if ((bomb_on == 1'b1) && (small_index != 0)) 
		begin
			Red = c_table[small_index][0];
			Green = c_table[small_index][1];
			Blue = c_table[small_index][2];
		end
		else if ((wall_on == 1'b1) && (big_index != 0)) 
		begin
			Red = c_table[big_index][0];
			Green = c_table[big_index][1];
			Blue = c_table[big_index][2];
		end
		else if ((tree_on == 1'b1) && (big_index != 0)) 
		begin
			Red = c_table[big_index][0];
			Green = c_table[big_index][1];
			Blue = c_table[big_index][2];
		end
		else if ((flame_on == 1'b1) && (small_index != 0)) 
		begin
			Red = c_table[small_index][0];
			Green = c_table[small_index][1];
			Blue = c_table[small_index][2];
		end
		else if ((coin_on == 1'b1) && (small_index != 0)) 
		begin
			Red = c_table[small_index][0];
			Green = c_table[small_index][1];
			Blue = c_table[small_index][2];
		end
		else if((score_on[0])&&(sprite_data[8-score_x_1]))
		begin
			Red = 8'd255;
			Green = 8'd223;
			Blue = 8'd0;
		end
		else if((score_on[1])&&(sprite_data[8-score_x_0]))
		begin
			Red = 8'd255;
			Green = 8'd223;
			Blue = 8'd0;
		end
		else if((score_on[2])&&(sprite_data[8-score_x_1]))
		begin
			Red = 8'd51;
			Green = 8'd255;
			Blue = 8'd255;
		end
		else if((score_on[3])&&(sprite_data[8-score_x_0]))
		begin
			Red = 8'd51;
			Green = 8'd255;
			Blue = 8'd255;
		end
		else if((coin_on)&&(sprite_data[8-((t1-12)/2)]))
		begin
			Red = 8'd225;
			Green = 8'd215;
			Blue = 8'd0;
		end
		else if((state == 2'b01)&&(Draw_X < 480))
		begin
			Red = c_table[tile_index][0];
			Green = c_table[tile_index][1];
			Blue = c_table[tile_index][2];
		end
		else if((player1_on)&&(~Player_choose)&&(sprite_scene[98-Draw_X + 272]))
		begin
			Red = 8'd255;
			Green = 8'd223;
			Blue = 8'd0;	
		end
		else if((player1_on)&&(Player_choose)&&(sprite_scene[98-Draw_X + 272]))
		begin
			Red = 8'd204;
			Green = 8'd206;
			Blue = 8'd143;	
		end
		else if((player2_on)&&(~Player_choose)&&(sprite_scene[98-Draw_X + 272]))
		begin
			Red = 8'd204;
			Green = 8'd206;
			Blue = 8'd143;	
		end
		else if((player2_on)&&(Player_choose)&&(sprite_scene[98-Draw_X + 272]))
		begin
			Red = 8'd255;
			Green = 8'd223;
			Blue = 8'd0;	
		end
		else if((final_on)&&(sprite_scene[98-(win_x/2)])&&(~Winner))
		begin
			Red = 8'd255;
			Green = 8'd223;
			Blue = 8'd0;	
		end
	   else if((final_on)&&(sprite_scene[98-(win_x/2)])&&(Winner))
		begin
			Red = 8'd51;
			Green = 8'd255;
			Blue = 8'd255;	
		end	
		else if((again_on)&&(sprite_2[98-again_x])&&(~Winner))
		begin
			Red = 8'd255;
			Green = 8'd223;
			Blue = 8'd0;	
		end
	   else if((again_on)&&(sprite_2[98-again_x])&&(Winner))
		begin
			Red = 8'd51;
			Green = 8'd255;
			Blue = 8'd255;	
		end	
		else
		begin
			Red = 8'd52;
			Green = 8'd61;
			Blue = 8'd70;
		end
	end 

endmodule
