module background(output logic [9:0] rgb[0:639][0:479]);
assign rgb = '{
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd426,9'd427,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd432,9'd433,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd434,9'd435,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd436,9'd437,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd438,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd439,9'd440,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd441,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd442,9'd443,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd444,9'd445,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd446,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd447,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd434,9'd443,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd448,9'd449,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd450,9'd445,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd444,9'd451,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd452,9'd453,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd436,9'd454,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd436,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd455,9'd456,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd444,9'd453,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd457,9'd458,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd459,9'd460,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd461,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd462,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd463,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd464,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd465,9'd466,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd467,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd468,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd469,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd448,9'd470,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd471,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd472,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd473,9'd470,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd474,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd452,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd467,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd475,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd477,9'd478,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd479,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd480,9'd453,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd481,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd482,9'd483,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd484,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd485,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd472,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd486,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd444,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd488,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd489,9'd483,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd490,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd491,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd492,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd493,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd494,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd427,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd495,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd463,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd461,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd434,9'd496,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd439,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd426,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd497,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd440,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd466,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd498,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd499,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd475,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd500,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd501,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd502,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd503,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd504,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd451,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd483,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd456,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd454,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd454,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd456,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd483,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd451,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd504,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd503,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd502,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd501,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd500,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd475,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd499,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd498,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd466,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd440,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd497,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd426,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd439,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd434,9'd496,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd461,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd463,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd495,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd427,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd494,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd493,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd492,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd491,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd490,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd489,9'd483,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd488,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd444,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd486,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd472,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd485,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd484,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd482,9'd483,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd481,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd480,9'd453,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd479,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd477,9'd478,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd475,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd467,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd452,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd474,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd473,9'd470,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd472,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd471,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd448,9'd470,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd469,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd468,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd467,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd465,9'd466,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd464,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd463,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd462,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd461,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd459,9'd460,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd457,9'd458,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd444,9'd453,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd455,9'd456,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd436,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd436,9'd454,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd452,9'd453,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd444,9'd451,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd450,9'd445,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd448,9'd449,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd434,9'd443,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd447,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd446,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd444,9'd445,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd442,9'd443,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd441,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd439,9'd440,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd438,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd436,9'd437,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd434,9'd435,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd432,9'd433,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd426,9'd427,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd428,9'd428,9'd428,9'd428,9'd428,9'd487,9'd487,9'd487,9'd487,9'd487,9'd487,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd476,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
},
'{
9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd425,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd429,9'd430,9'd430,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431,9'd431
}};
endmodule
