module Color_Table (
	output logic [7:0] colors[0:8][0:2]
);

assign colors = '{'{8'd255,8'd0,8'd0},'{8'd0,8'd26,8'd0},'{8'd241,8'd241,8'd231},'{8'd226,8'd133,8'd77},'{8'd226,8'd133,8'd77},
'{8'd73,8'd73,8'd36}, '{8'd225,8'd223,8'd0}, '{8'd225,8'd223,8'd0}, '{8'd61,8'd86,8'd52}};


endmodule
