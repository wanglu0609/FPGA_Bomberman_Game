module bird_sprite2(output logic [9:0] rgb[0:31][0:31]);
assign rgb = '{
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd254,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd255,9'd5,9'd256,9'd256,9'd257,9'd8,9'd258,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd259,9'd259,9'd260,9'd261,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd258,9'd262,9'd256,9'd263,9'd264,9'd265,9'd266,9'd256,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd18,9'd267,9'd18,9'd268,9'd21,9'd21,9'd22,9'd21,9'd261,9'd261,9'd260,9'd5,9'd5,9'd269,9'd270,9'd271,9'd28,9'd26,9'd28,9'd272,9'd273,9'd8,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd33,9'd274,9'd24,9'd24,9'd275,9'd276,9'd37,9'd260,9'd260,9'd268,9'd267,9'd269,9'd5,9'd269,9'd277,9'd278,9'd279,9'd26,9'd26,9'd26,9'd264,9'd280,9'd5,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd18,9'd260,9'd47,9'd37,9'd281,9'd281,9'd276,9'd48,9'd37,9'd260,9'd282,9'd262,9'd256,9'd283,9'd265,9'd28,9'd26,9'd26,9'd26,9'd26,9'd26,9'd279,9'd284,9'd256,9'd5,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd281,9'd22,9'd22,9'd22,9'd22,9'd260,9'd53,9'd285,9'd53,9'd37,9'd261,9'd261,9'd286,9'd287,9'd288,9'd26,9'd26,9'd26,9'd26,9'd26,9'd26,9'd279,9'd289,9'd290,9'd291,9'd273,9'd292
},
'{
9'd0,9'd0,9'd0,9'd0,9'd267,9'd58,9'd58,9'd22,9'd59,9'd60,9'd61,9'd62,9'd53,9'd293,9'd48,9'd37,9'd140,9'd294,9'd288,9'd26,9'd26,9'd26,9'd26,9'd26,9'd26,9'd26,9'd295,9'd43,9'd43,9'd296,9'd297,9'd0
},
'{
9'd0,9'd0,9'd0,9'd274,9'd22,9'd58,9'd59,9'd70,9'd298,9'd72,9'd73,9'd72,9'd299,9'd74,9'd53,9'd294,9'd262,9'd273,9'd287,9'd28,9'd26,9'd26,9'd26,9'd26,9'd26,9'd28,9'd28,9'd300,9'd301,9'd302,9'd0,9'd0
},
'{
9'd0,9'd0,9'd79,9'd58,9'd58,9'd70,9'd22,9'd81,9'd82,9'd83,9'd84,9'd83,9'd85,9'd303,9'd87,9'd304,9'd305,9'd280,9'd306,9'd279,9'd26,9'd26,9'd26,9'd26,9'd26,9'd26,9'd26,9'd307,9'd293,9'd5,9'd308,9'd0
},
'{
9'd0,9'd89,9'd275,9'd21,9'd261,9'd70,9'd22,9'd90,9'd91,9'd309,9'd93,9'd93,9'd84,9'd94,9'd310,9'd311,9'd312,9'd313,9'd28,9'd26,9'd26,9'd279,9'd26,9'd279,9'd28,9'd295,9'd314,9'd43,9'd315,9'd297,9'd0,9'd0
},
'{
9'd0,9'd316,9'd268,9'd261,9'd260,9'd260,9'd58,9'd317,9'd318,9'd102,9'd103,9'd104,9'd93,9'd83,9'd85,9'd319,9'd5,9'd320,9'd28,9'd321,9'd322,9'd28,9'd28,9'd323,9'd324,9'd43,9'd43,9'd44,9'd325,9'd326,9'd261,9'd0
},
'{
9'd0,9'd327,9'd47,9'd268,9'd37,9'd70,9'd58,9'd328,9'd112,9'd113,9'd114,9'd115,9'd116,9'd329,9'd330,9'd331,9'd5,9'd270,9'd332,9'd43,9'd43,9'd333,9'd321,9'd334,9'd43,9'd43,9'd334,9'd335,9'd280,9'd266,9'd260,9'd0
},
'{
9'd47,9'd283,9'd37,9'd336,9'd53,9'd70,9'd59,9'd125,9'd337,9'd127,9'd128,9'd338,9'd339,9'd340,9'd132,9'd341,9'd342,9'd5,9'd343,9'd44,9'd314,9'd344,9'd44,9'd43,9'd44,9'd296,9'd292,9'd269,9'd256,9'd17,9'd345,9'd0
},
'{
9'd37,9'd24,9'd75,9'd48,9'd53,9'd140,9'd74,9'd141,9'd142,9'd127,9'd113,9'd128,9'd143,9'd143,9'd144,9'd141,9'd346,9'd283,9'd270,9'd344,9'd269,9'd256,9'd315,9'd301,9'd347,9'd348,9'd269,9'd269,9'd0,9'd0,9'd0,9'd0
},
'{
9'd47,9'd349,9'd17,9'd275,9'd53,9'd48,9'd74,9'd150,9'd132,9'd337,9'd127,9'd350,9'd152,9'd337,9'd153,9'd351,9'd352,9'd353,9'd354,9'd338,9'd291,9'd262,9'd355,9'd356,9'd256,9'd5,9'd356,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd70,9'd79,9'd308,9'd24,9'd285,9'd159,9'd60,9'd160,9'd357,9'd162,9'd358,9'd163,9'd164,9'd102,9'd359,9'd360,9'd163,9'd361,9'd358,9'd157,9'd362,9'd346,9'd362,9'd329,9'd283,9'd363,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd336,9'd364,9'd308,9'd5,9'd17,9'd17,9'd17,9'd62,9'd365,9'd162,9'd350,9'd358,9'd173,9'd174,9'd175,9'd128,9'd163,9'd358,9'd350,9'd366,9'd218,9'd318,9'd367,9'd368,9'd328,9'd319,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd140,9'd18,9'd283,9'd308,9'd283,9'd293,9'd17,9'd159,9'd179,9'd369,9'd350,9'd114,9'd157,9'd370,9'd181,9'd115,9'd182,9'd114,9'd173,9'd174,9'd183,9'd371,9'd370,9'd368,9'd346,9'd317,9'd372,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd260,9'd349,9'd348,9'd283,9'd373,9'd293,9'd159,9'd189,9'd190,9'd191,9'd192,9'd370,9'd193,9'd192,9'd115,9'd194,9'd194,9'd195,9'd196,9'd197,9'd365,9'd193,9'd199,9'd374,9'd85,9'd372,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd21,9'd276,9'd275,9'd280,9'd375,9'd373,9'd75,9'd189,9'd160,9'd203,9'd103,9'd352,9'd102,9'd337,9'd173,9'd194,9'd157,9'd204,9'd352,9'd205,9'd205,9'd206,9'd338,9'd367,9'd207,9'd208,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd47,9'd260,9'd276,9'd75,9'd5,9'd272,9'd285,9'd140,9'd210,9'd82,9'd299,9'd360,9'd212,9'd213,9'd337,9'd173,9'd352,9'd215,9'd376,9'd152,9'd377,9'd217,9'd164,9'd218,9'd378,9'd303,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd58,9'd276,9'd379,9'd75,9'd17,9'd159,9'd60,9'd219,9'd219,9'd220,9'd380,9'd358,9'd213,9'd173,9'd361,9'd222,9'd381,9'd382,9'd278,9'd225,9'd382,9'd222,9'd338,9'd383,9'd384,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd22,9'd37,9'd379,9'd140,9'd17,9'd60,9'd60,9'd219,9'd228,9'd229,9'd361,9'd366,9'd114,9'd385,9'd230,9'd231,9'd232,9'd233,9'd234,9'd386,9'd339,9'd338,9'd183,9'd319,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd276,9'd261,9'd37,9'd70,9'd140,9'd189,9'd74,9'd74,9'd179,9'd387,9'd350,9'd163,9'd174,9'd173,9'd191,9'd357,9'd237,9'd238,9'd237,9'd239,9'd157,9'd366,9'd388,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd47,9'd58,9'd260,9'd70,9'd70,9'd59,9'd240,9'd219,9'd72,9'd191,9'd241,9'd352,9'd380,9'd197,9'd242,9'd243,9'd244,9'd239,9'd241,9'd245,9'd128,9'd203,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd58,9'd261,9'd58,9'd58,9'd261,9'd22,9'd74,9'd22,9'd303,9'd371,9'd371,9'd318,9'd112,9'd128,9'd369,9'd164,9'd218,9'd182,9'd157,9'd229,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd260,9'd22,9'd22,9'd22,9'd58,9'd22,9'd74,9'd247,9'd70,9'd248,9'd389,9'd389,9'd362,9'd362,9'd383,9'd252,9'd252,9'd383,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd47,9'd22,9'd58,9'd22,9'd58,9'd58,9'd22,9'd247,9'd247,9'd247,9'd253,9'd48,9'd390,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd260,9'd22,9'd22,9'd22,9'd22,9'd140,9'd260,9'd22,9'd247,9'd22,9'd22,9'd22,9'd22,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd58,9'd22,9'd22,9'd336,9'd276,9'd260,9'd22,9'd58,9'd261,9'd261,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
},
'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd261,9'd261,9'd0,9'd0,9'd260,9'd47,9'd47,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0
}};
endmodule
