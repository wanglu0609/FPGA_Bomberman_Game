module exploded (output logic [7:0] index[0:39][0:39]);

assign index = '{
'{
8'd21,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd21,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd21,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd21,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd22,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd21,8'd21,8'd21,8'd21,8'd21,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd21,8'd23,8'd23,8'd23,8'd23,8'd23,8'd23,8'd21,8'd21,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd23,8'd23,8'd21,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd23,8'd21,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd4,8'd4,8'd4,8'd4,8'd18,8'd18,8'd23,8'd21,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd4,8'd4,8'd4,8'd4,8'd4,8'd4,8'd18,8'd23,8'd21,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd4,8'd4,8'd4,8'd4,8'd4,8'd4,8'd18,8'd18,8'd23,8'd21,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd4,8'd4,8'd4,8'd4,8'd4,8'd4,8'd18,8'd18,8'd23,8'd21,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd22,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd4,8'd4,8'd4,8'd4,8'd4,8'd4,8'd18,8'd18,8'd23,8'd21,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd22,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd4,8'd4,8'd4,8'd4,8'd18,8'd18,8'd18,8'd23,8'd21,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd23,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd23,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd23,8'd21,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd23,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd23,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd18,8'd18,8'd18,8'd18,8'd18,8'd18,8'd23,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd23,8'd23,8'd23,8'd23,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd22,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd22,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd19,8'd22,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd19,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd22,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd22,8'd22,8'd22},

'{
8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd19,8'd22,8'd22},

'{
8'd20,8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd19,8'd22},

'{
8'd20,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd22},

'{
8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21,8'd21}
};

endmodule
