module Char_Sprite(
	output logic [8:0] index[0:47][0:47]
);

assign index = '{

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd3,9'd3,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd3,9'd3,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd3,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd3,9'd6,9'd3,9'd3,9'd6,9'd6,9'd6,9'd6,9'd3,9'd3,9'd6,9'd3,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd6,9'd6,9'd3,9'd3,9'd6,9'd6,9'd6,9'd6,9'd3,9'd3,9'd6,9'd6,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd6,9'd6,9'd3,9'd3,9'd6,9'd6,9'd6,9'd6,9'd3,9'd3,9'd6,9'd6,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd3,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd6,9'd3,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd0,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd2,9'd0,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd2,9'd2,9'd2,9'd0,9'd0,9'd2,9'd2,9'd2,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd8,9'd2,9'd2,9'd2,9'd3,9'd8,9'd2,9'd2,9'd2,9'd3,9'd8,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd8,9'd8,9'd2,9'd2,9'd2,9'd8,9'd8,9'd2,9'd2,9'd2,9'd8,9'd8,9'd8,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd8,9'd8,9'd3,9'd3,9'd8,9'd8,9'd8,9'd3,9'd3,9'd8,9'd8,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0},

'{
9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0,9'd0}


};

endmodule
