module color_table (output logic [7:0] colors[0:33][0:2]);

assign colors = '{'{8'd255,8'd0,8'd0},
'{8'd41, 8'd37, 8'd37},
'{8'd75, 8'd70, 8'd70},
'{8'd255, 8'd223, 8'd0},
'{8'd215, 8'd93, 8'd0},
'{8'd228, 8'd151, 8'd97},
'{8'd249, 8'd249, 8'd238},
'{8'd228, 8'd226, 8'd192},
'{8'd63, 8'd88, 8'd55},
'{8'd60, 8'd109, 8'd72},
'{8'd71, 8'd122, 8'd82},
'{8'd20, 8'd18, 8'd40},
'{8'd44, 8'd43, 8'd70},
'{8'd30, 8'd28, 8'd51},
'{8'd63, 8'd63, 8'd87},
'{8'd16, 8'd15, 8'd37},
'{8'd11, 8'd8, 8'd31},
'{8'd215, 8'd93, 8'd0},
'{8'd173, 8'd78, 8'd6},
'{8'd104, 8'd127, 8'd144},
'{8'd79, 8'd94, 8'd105},
'{8'd85, 8'd107, 8'd123},
'{8'd112, 8'd132, 8'd147},
'{8'd99, 8'd103, 8'd111},
'{8'd209, 8'd0, 8'd0},
'{8'd255, 8'd206, 8'd0},
'{8'd217, 8'd60, 8'd0},
'{8'd255, 8'd191, 8'd0},
'{8'd255, 8'd209, 8'd0},
'{8'd146, 8'd73, 8'd0},
'{8'd20, 8'd18, 8'd40},
'{8'd255, 8'd255, 8'd255},
'{8'd228, 8'd226, 8'd192},
'{8'd57, 8'd37, 8'd129}};


endmodule
