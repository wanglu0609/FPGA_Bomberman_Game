module five(output logic [9:0] rgb[0:23][0:31]);
assign rgb = '{
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd428,9'd430,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd428,9'd428,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd428,9'd428,9'd430,9'd430,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd428,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd428,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd428,9'd428,9'd428,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd430,9'd430,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd430,9'd428,9'd428,9'd428,9'd428,9'd428,9'd428,9'd430,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd430,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
}};
endmodule
