module flame (output logic [7:0] index[0:27][0:27]);

assign index = '{
'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd26,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd4,8'd26,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd26,8'd26,8'd26,8'd26,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd25,8'd25,8'd0,8'd0,8'd26,8'd26,8'd26,8'd26,8'd26,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd28,8'd28,8'd25,8'd0,8'd26,8'd26,8'd26,8'd26,8'd26,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd29,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd24,8'd0,8'd0,8'd3,8'd25,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd0,8'd0,8'd18,8'd18,8'd29,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd24,8'd26,8'd28,8'd27,8'd4,8'd26,8'd26,8'd26,8'd26,8'd4,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd29,8'd18,8'd29,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd24,8'd24,8'd27,8'd25,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd4,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd18,8'd18,8'd29,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd24,8'd26,8'd27,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd27,8'd27,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd18,8'd18,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd24,8'd4,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd4,8'd28,8'd25,8'd4,8'd26,8'd4,8'd26,8'd26,8'd26,8'd26,8'd18,8'd24,8'd24,8'd24,8'd0},

'{
8'd0,8'd0,8'd0,8'd24,8'd24,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd4,8'd25,8'd25,8'd25,8'd27,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd24,8'd24,8'd0},

'{
8'd0,8'd0,8'd0,8'd24,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd4,8'd25,8'd25,8'd25,8'd25,8'd28,8'd27,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd24,8'd24,8'd0},

'{
8'd0,8'd0,8'd24,8'd24,8'd26,8'd26,8'd26,8'd26,8'd26,8'd26,8'd4,8'd25,8'd25,8'd25,8'd25,8'd25,8'd25,8'd28,8'd27,8'd4,8'd26,8'd26,8'd26,8'd26,8'd4,8'd26,8'd24,8'd24},

'{
8'd0,8'd24,8'd24,8'd26,8'd4,8'd26,8'd26,8'd26,8'd26,8'd4,8'd25,8'd25,8'd25,8'd25,8'd28,8'd25,8'd25,8'd25,8'd25,8'd27,8'd4,8'd26,8'd26,8'd26,8'd26,8'd26,8'd24,8'd24},

'{
8'd0,8'd24,8'd24,8'd26,8'd26,8'd26,8'd26,8'd26,8'd4,8'd25,8'd25,8'd25,8'd25,8'd28,8'd3,8'd28,8'd25,8'd25,8'd25,8'd28,8'd27,8'd4,8'd26,8'd26,8'd26,8'd4,8'd26,8'd24},

'{
8'd0,8'd24,8'd24,8'd26,8'd26,8'd26,8'd26,8'd4,8'd25,8'd25,8'd25,8'd25,8'd28,8'd3,8'd3,8'd3,8'd28,8'd25,8'd25,8'd25,8'd28,8'd27,8'd26,8'd26,8'd26,8'd4,8'd26,8'd0},

'{
8'd24,8'd24,8'd24,8'd26,8'd26,8'd26,8'd26,8'd27,8'd28,8'd25,8'd25,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd28,8'd25,8'd25,8'd25,8'd28,8'd4,8'd26,8'd26,8'd4,8'd26,8'd0},

'{
8'd24,8'd24,8'd24,8'd26,8'd4,8'd26,8'd4,8'd25,8'd25,8'd25,8'd25,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd25,8'd25,8'd25,8'd28,8'd27,8'd26,8'd26,8'd4,8'd0,8'd0},

'{
8'd24,8'd24,8'd24,8'd26,8'd4,8'd26,8'd4,8'd25,8'd25,8'd25,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd28,8'd25,8'd25,8'd28,8'd27,8'd26,8'd26,8'd4,8'd0,8'd0},

'{
8'd0,8'd24,8'd24,8'd24,8'd26,8'd26,8'd4,8'd25,8'd25,8'd25,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd28,8'd25,8'd25,8'd28,8'd27,8'd26,8'd26,8'd26,8'd0,8'd0},

'{
8'd0,8'd24,8'd24,8'd24,8'd26,8'd4,8'd26,8'd27,8'd25,8'd25,8'd25,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd25,8'd25,8'd25,8'd28,8'd27,8'd26,8'd4,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd24,8'd24,8'd24,8'd26,8'd26,8'd4,8'd28,8'd25,8'd25,8'd25,8'd28,8'd3,8'd3,8'd3,8'd28,8'd25,8'd25,8'd25,8'd25,8'd28,8'd4,8'd26,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd24,8'd24,8'd24,8'd26,8'd4,8'd27,8'd28,8'd25,8'd25,8'd25,8'd25,8'd25,8'd25,8'd25,8'd25,8'd25,8'd28,8'd28,8'd27,8'd26,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd24,8'd24,8'd24,8'd26,8'd4,8'd27,8'd28,8'd28,8'd25,8'd25,8'd25,8'd25,8'd25,8'd28,8'd28,8'd27,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd27,8'd27,8'd27,8'd27,8'd27,8'd27,8'd27,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0}


};

endmodule
