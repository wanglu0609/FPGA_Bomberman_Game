module tile (output logic [7:0] index[0:39][0:39]);

assign index = '{
'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd9,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd9,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd9,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd9,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd9,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10},

'{
8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10,8'd10}

};

endmodule
