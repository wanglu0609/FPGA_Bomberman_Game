module bomb_sprites (output logic [7:0] index[0:27][0:27]);

assign index = '{
'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd15,8'd15,8'd15,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd13,8'd13,8'd13,8'd11,8'd15,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd11,8'd15,8'd16,8'd16,8'd12,8'd33,8'd33,8'd33,8'd33,8'd13,8'd15,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd15,8'd13,8'd22,8'd22,8'd21,8'd33,8'd33,8'd33,8'd33,8'd33,8'd13,8'd15,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd11,8'd11,8'd7,8'd7,8'd7,8'd7,8'd22,8'd33,8'd33,8'd33,8'd33,8'd14,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0},

'{
8'd0,8'd11,8'd16,8'd2,8'd7,8'd20,8'd33,8'd21,8'd7,8'd22,8'd33,8'd33,8'd33,8'd33,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0},

'{
8'd0,8'd11,8'd16,8'd20,8'd7,8'd21,8'd33,8'd33,8'd22,8'd22,8'd33,8'd33,8'd33,8'd33,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0},

'{
8'd0,8'd11,8'd11,8'd13,8'd7,8'd22,8'd33,8'd33,8'd33,8'd33,8'd33,8'd33,8'd33,8'd33,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0},

'{
8'd0,8'd11,8'd11,8'd16,8'd20,8'd7,8'd33,8'd33,8'd33,8'd33,8'd33,8'd33,8'd33,8'd13,8'd15,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0},

'{
8'd11,8'd11,8'd15,8'd23,8'd7,8'd7,8'd14,8'd33,8'd33,8'd33,8'd33,8'd33,8'd12,8'd15,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11},

'{
8'd11,8'd15,8'd12,8'd31,8'd31,8'd7,8'd15,8'd11,8'd13,8'd12,8'd12,8'd13,8'd15,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11},

'{
8'd11,8'd15,8'd11,8'd7,8'd31,8'd22,8'd16,8'd11,8'd15,8'd15,8'd15,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11},

'{
8'd11,8'd11,8'd15,8'd13,8'd14,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11},

'{
8'd0,8'd11,8'd11,8'd15,8'd16,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0},

'{
8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0},

'{
8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0},

'{
8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0},

'{
8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd11,8'd11,8'd11,8'd11,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0}


};

endmodule
