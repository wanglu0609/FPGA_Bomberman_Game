module right (output logic [7:0] index[0:179][0:39]);

assign index = '{'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd7,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd4,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd5,8'd26,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd5,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd28,8'd5,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd25,8'd23,8'd25,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd5,8'd21,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd5,8'd21,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd25,8'd23,8'd25,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd5,8'd3,8'd3,8'd3,8'd28,8'd5,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd5,8'd3,8'd3,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd7,8'd7,8'd7,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd7,8'd7,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd15,8'd22,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd31,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd1,8'd22,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd7,8'd23,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd1,8'd22,8'd7,8'd7,8'd7,8'd7,8'd7,8'd22,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd10,8'd7,8'd7,8'd7,8'd7,8'd5,8'd1,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd23,8'd7,8'd7,8'd22,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd1,8'd1,8'd1,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd7,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd4,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd5,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd28,8'd28,8'd28,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd28,8'd5,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd5,8'd21,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd5,8'd21,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd5,8'd21,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd28,8'd22,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd28,8'd3,8'd3,8'd3,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd1,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd10,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd1,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd10,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd1,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd9,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd1,8'd22,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd22,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd7,8'd6,8'd31,8'd6,8'd7,8'd7,8'd22,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd22,8'd22,8'd23,8'd1,8'd1,8'd1,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd1,8'd15,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd7,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd4,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd5,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd4,8'd4,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd28,8'd28,8'd28,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd28,8'd5,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd5,8'd21,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd5,8'd21,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd5,8'd21,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd28,8'd22,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd28,8'd3,8'd3,8'd3,8'd28,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd5,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd3,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd31,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd31,8'd31,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd7,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd31,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd22,8'd6,8'd6,8'd6,8'd6,8'd6,8'd7,8'd7,8'd7,8'd7,8'd7,8'd22,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd22,8'd6,8'd6,8'd6,8'd6,8'd6,8'd22,8'd10,8'd7,8'd7,8'd22,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd23,8'd6,8'd6,8'd6,8'd6,8'd6,8'd22,8'd16,8'd1,8'd1,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd7,8'd31,8'd6,8'd6,8'd31,8'd22,8'd1,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd1,8'd22,8'd6,8'd31,8'd6,8'd7,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd8,8'd8,8'd1,8'd23,8'd22,8'd22,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd8,8'd8,8'd8,8'd16,8'd1,8'd8,8'd8,8'd8,8'd8,8'd8,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0},

'{
8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0,8'd0}




};

endmodule
