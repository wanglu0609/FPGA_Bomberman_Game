module fireball(output logic [9:0] rgb[0:31][0:31]);
assign rgb = '{
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd392,9'd392,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd393,9'd393,9'd391,9'd391,9'd393,9'd394,9'd393,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd393,9'd391,9'd391,9'd391,9'd392,9'd394,9'd394,9'd394,9'd393,9'd392,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd393,9'd393,9'd392,9'd392,9'd393,9'd393,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd393,9'd393,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd393,9'd394,9'd394,9'd393,9'd393,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd395,9'd395,9'd395,9'd395,9'd394,9'd394,9'd393,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd396,9'd396,9'd396,9'd395,9'd395,9'd395,9'd394,9'd394,9'd393,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd393,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd395,9'd396,9'd397,9'd397,9'd396,9'd396,9'd396,9'd395,9'd394,9'd394,9'd393,9'd392,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd393,9'd394,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd395,9'd395,9'd396,9'd396,9'd397,9'd397,9'd396,9'd396,9'd396,9'd395,9'd395,9'd394,9'd394,9'd393,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd395,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd396,9'd396,9'd396,9'd396,9'd396,9'd397,9'd397,9'd397,9'd397,9'd396,9'd396,9'd395,9'd394,9'd394,9'd393,9'd392,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd392,9'd391,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd396,9'd396,9'd397,9'd397,9'd396,9'd396,9'd397,9'd397,9'd136,9'd136,9'd397,9'd396,9'd395,9'd394,9'd394,9'd394,9'd394,9'd393,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd392,9'd392,9'd392,9'd394,9'd394,9'd394,9'd395,9'd395,9'd395,9'd396,9'd397,9'd397,9'd397,9'd396,9'd396,9'd397,9'd397,9'd397,9'd136,9'd397,9'd396,9'd396,9'd395,9'd394,9'd394,9'd394,9'd395,9'd392,9'd391
},
'{
9'd391,9'd391,9'd391,9'd393,9'd392,9'd393,9'd395,9'd394,9'd394,9'd395,9'd395,9'd396,9'd396,9'd397,9'd397,9'd397,9'd397,9'd136,9'd136,9'd397,9'd397,9'd396,9'd396,9'd136,9'd396,9'd396,9'd395,9'd394,9'd394,9'd394,9'd393,9'd391
},
'{
9'd391,9'd391,9'd393,9'd394,9'd393,9'd394,9'd395,9'd395,9'd395,9'd395,9'd395,9'd396,9'd397,9'd397,9'd136,9'd136,9'd398,9'd399,9'd399,9'd398,9'd397,9'd396,9'd396,9'd397,9'd396,9'd396,9'd396,9'd395,9'd394,9'd394,9'd394,9'd391
},
'{
9'd391,9'd391,9'd393,9'd394,9'd394,9'd394,9'd395,9'd396,9'd396,9'd396,9'd395,9'd396,9'd397,9'd397,9'd136,9'd398,9'd398,9'd399,9'd399,9'd398,9'd397,9'd396,9'd396,9'd397,9'd397,9'd396,9'd396,9'd395,9'd394,9'd394,9'd394,9'd393
},
'{
9'd391,9'd391,9'd394,9'd394,9'd394,9'd394,9'd395,9'd396,9'd397,9'd396,9'd396,9'd396,9'd397,9'd397,9'd398,9'd398,9'd399,9'd399,9'd399,9'd136,9'd397,9'd397,9'd397,9'd397,9'd397,9'd397,9'd396,9'd396,9'd395,9'd394,9'd394,9'd393
},
'{
9'd391,9'd392,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd396,9'd396,9'd396,9'd397,9'd397,9'd398,9'd399,9'd399,9'd399,9'd399,9'd399,9'd136,9'd397,9'd136,9'd136,9'd397,9'd397,9'd397,9'd396,9'd396,9'd395,9'd394,9'd394,9'd393
},
'{
9'd391,9'd393,9'd394,9'd394,9'd394,9'd394,9'd394,9'd395,9'd396,9'd396,9'd397,9'd397,9'd398,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd136,9'd397,9'd397,9'd396,9'd396,9'd395,9'd394,9'd394,9'd393
},
'{
9'd391,9'd393,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd395,9'd396,9'd396,9'd397,9'd136,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd136,9'd397,9'd397,9'd396,9'd396,9'd395,9'd394,9'd394,9'd393
},
'{
9'd391,9'd391,9'd394,9'd394,9'd395,9'd395,9'd395,9'd395,9'd396,9'd396,9'd396,9'd397,9'd136,9'd398,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd398,9'd397,9'd397,9'd396,9'd397,9'd396,9'd395,9'd394,9'd394,9'd391
},
'{
9'd391,9'd391,9'd393,9'd394,9'd395,9'd395,9'd395,9'd396,9'd396,9'd396,9'd396,9'd396,9'd397,9'd136,9'd398,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd399,9'd136,9'd397,9'd397,9'd396,9'd397,9'd397,9'd395,9'd394,9'd393,9'd391
},
'{
9'd391,9'd391,9'd393,9'd395,9'd395,9'd396,9'd397,9'd396,9'd396,9'd396,9'd396,9'd396,9'd396,9'd397,9'd136,9'd398,9'd398,9'd399,9'd399,9'd399,9'd399,9'd399,9'd136,9'd397,9'd396,9'd396,9'd396,9'd396,9'd394,9'd394,9'd393,9'd391
},
'{
9'd391,9'd391,9'd392,9'd395,9'd396,9'd396,9'd397,9'd136,9'd397,9'd396,9'd396,9'd396,9'd395,9'd395,9'd396,9'd397,9'd397,9'd136,9'd398,9'd399,9'd399,9'd398,9'd136,9'd397,9'd396,9'd395,9'd396,9'd396,9'd394,9'd394,9'd391,9'd391
},
'{
9'd391,9'd391,9'd392,9'd393,9'd395,9'd396,9'd396,9'd397,9'd396,9'd396,9'd395,9'd395,9'd395,9'd395,9'd395,9'd396,9'd397,9'd397,9'd136,9'd136,9'd136,9'd136,9'd136,9'd396,9'd396,9'd396,9'd396,9'd395,9'd394,9'd393,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd393,9'd394,9'd395,9'd395,9'd395,9'd395,9'd395,9'd395,9'd395,9'd396,9'd396,9'd396,9'd397,9'd397,9'd397,9'd397,9'd397,9'd397,9'd397,9'd397,9'd396,9'd395,9'd396,9'd396,9'd394,9'd394,9'd393,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd392,9'd393,9'd393,9'd394,9'd394,9'd394,9'd395,9'd395,9'd395,9'd396,9'd396,9'd397,9'd397,9'd397,9'd397,9'd397,9'd397,9'd397,9'd396,9'd396,9'd395,9'd395,9'd393,9'd392,9'd393,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd393,9'd394,9'd394,9'd394,9'd395,9'd395,9'd395,9'd396,9'd396,9'd397,9'd397,9'd397,9'd397,9'd396,9'd396,9'd395,9'd395,9'd394,9'd392,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd392,9'd393,9'd394,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd396,9'd396,9'd397,9'd397,9'd396,9'd396,9'd395,9'd395,9'd394,9'd393,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd393,9'd394,9'd394,9'd394,9'd394,9'd394,9'd395,9'd395,9'd396,9'd396,9'd396,9'd396,9'd395,9'd394,9'd394,9'd394,9'd393,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd392,9'd393,9'd394,9'd394,9'd394,9'd395,9'd395,9'd395,9'd395,9'd395,9'd394,9'd394,9'd394,9'd393,9'd392,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd392,9'd393,9'd393,9'd394,9'd394,9'd394,9'd394,9'd394,9'd394,9'd393,9'd393,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd392,9'd393,9'd394,9'd393,9'd393,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
}};
endmodule
