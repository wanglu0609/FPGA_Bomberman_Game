module bottom_pipe(output logic [9:0] rgb[0:47][0:379]);
assign rgb = '{
'{
9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd400,9'd400,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd400,9'd400,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd400,9'd400,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400
},
'{
9'd400,9'd400,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd400,9'd400,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402,9'd402
},
'{
9'd400,9'd400,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd403,9'd400,9'd400,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404,9'd404
},
'{
9'd400,9'd400,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd400,9'd400,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401
},
'{
9'd400,9'd400,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd401,9'd400,9'd400,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405,9'd405
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407,9'd407
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408,9'd408
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409,9'd409
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410,9'd410
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411,9'd411
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412,9'd412
},
'{
9'd400,9'd400,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd406,9'd400,9'd400,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413,9'd413
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415,9'd415
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416,9'd416
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417,9'd417
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418,9'd418
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419,9'd419
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420,9'd420
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421
},
'{
9'd400,9'd400,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd400,9'd400,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421
},
'{
9'd400,9'd400,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd400,9'd400,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421,9'd421
},
'{
9'd400,9'd400,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd422,9'd400,9'd400,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423,9'd423
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424,9'd424
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400
},
'{
9'd400,9'd400,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd414,9'd400,9'd400,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
},
'{
9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd400,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391,9'd391
}};
endmodule
