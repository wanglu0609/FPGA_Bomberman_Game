module Solid (output logic [7:0] index[0:39][0:39]);

assign index = '{
'{
8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd15,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd15,8'd11,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd15,8'd11,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd15,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd11,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd13,8'd11,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd12,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd14,8'd13,8'd16,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd13,8'd15,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd13,8'd11,8'd11,8'd15,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd13,8'd16,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12,8'd12},

'{
8'd11,8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12,8'd12},

'{
8'd11,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd12},

'{
8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13,8'd13}
};
endmodule
